module cuMV(
    input logic                 clk,
    input logic                 RegWriteM,
    input logic     [1:0]       ResultSrcM,

    output logic                RegWriteW,
    output logic    [1:0]       ResultSrcW,
);

// do we create register for each signal since each have different width size?

endmodule
